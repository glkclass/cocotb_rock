// User lib. Add missed units here

// replace missed stuff
module BUF_X0_12_LVT_NT (input A, output Q);
	assign Q = A;
endmodule

